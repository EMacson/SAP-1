`timescale 1ns / 1ps

module d_latch (
    input d,
    output wire q,
    output wire q`
);

endmodule